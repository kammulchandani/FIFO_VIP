`include "../top/defines.sv"
`include "./fifo_seq_item.sv"
`include "./fifo_sequencer.sv"
`include "./fifo_vsequencer.sv"
`include "./fifo_driver.sv"
`include "./fifo_drvr_monitor.sv"
`include "./fifo_dut_monitor.sv"
`include "./fifo_drvr_agent.sv"
`include "./fifo_dut_agent.sv"
`include "./fifo_uvc.sv"
`include "./../top/fifo_sb.sv"
`include "./../top/fifo_tb.sv"
`include "./../sequences/fifo_seqs.sv"
`include "./../sequences/fifo_vseqs.sv"
